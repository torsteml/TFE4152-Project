//-----------------------------------------------------------------------------
//
// Title       : Timer_counter
// Design      : camera
// Author      : markusru
// Company     : NTNU
//
//-----------------------------------------------------------------------------
//
// File        : c:\My_Designs\ICprosjekt\camera\src\Timer_counter.v
// Generated   : Tue Nov  6 15:13:38 2018
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {Timer_counter}}
module Timer_counter ( Reset ,clk ,Start ,Initial ,Ovf5 );

output Ovf5 ;
wire Ovf5 ;

input Reset ;
wire Reset ;
input clk ;
wire clk ;
input Start ;
wire Start ;
input Initial ;
wire Initial ;

//}} End of automatically maintained section

// -- Enter your statements here -- //

begin @(Start)


	
end

endmodule
