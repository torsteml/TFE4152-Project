[aimspice]
[description]
2053
Analog part

.include p18_cmos_models_tt.inc
.include p18_model_card.inc

X11 VDD 0 Expose Erase NRE_R1 OUT1 OnePixel
X12 VDD 0 Expose Erase NRE_R1 OUT2 OnePixel
X21 VDD 0 Expose Erase NRE_R2 OUT1 OnePixel
X22 VDD 0 Expose Erase NRE_R2 OUT2 OnePixel
XLT1 VDD 0 OUT1 LoadTransistor
XLT2 VDD 0 OUT2 LoadTransistor


.param Ipd_1 = 750p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 2m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_R1_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R1 signal
.param NRE_R2_DLY = {4*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE_R2 signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD VDD 0 dc VDD
VEXPOSE EXPOSE 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE ERASE 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R1 NRE_R1 0 dc 0 pulse(VDD 0 NRE_R1_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE_R2 NRE_R2 0 dc 0  pulse(VDD 0 NRE_R2_DLY TRF TRF CLK_PERIOD PERIOD)

.plot V(EXPOSE) V(NRE_R1) V(NRE_R2) V(ERASE)
.plot V(OUT1) V(OUT2) ! signals going to ADC
.plot V(OUT_SAMPLED1)

.subckt LoadTransistor Vdd Vss Gate
MC Gate Gate Vdd Vdd PMOS L=2u W=10u
CC Gate Vss 3p
.ends

.subckt OnePixel Vdd Vss Expose Erase NRE Out
XPD1 Vdd N1 PhotoDiode
MN1 N1 Expose N2 Vss NMOS L=0.7u W=10u
MN2 N2 Erase Vss Vss NMOS L=2u W=2u
CS N2 Vss 0.833p
MP3 Vss N2 N3 Vdd PMOS L=2u W=10u
MP4 N3 NRE Out Vdd PMOS L=0.7u W=10u
.ends

.subckt PhotoDiode  VDD N1_R1C1
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends 



[dc]
1
VDD
1
2
0.1
[tran]
0.0001
0.060
X
X
0
[ana]
4 0
[end]
