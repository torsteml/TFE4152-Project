[aimspice]
[description]
1483
OnePixel

.include p18_cmos_models_tt.inc
.include p18_model_card.inc

XPD1 Vdd N1 PhotoDiode
MN1 N1 Expose N2 0 NMOS L=0.7u W=10u
MN2 N2 Erase 0 0 NMOS L=2u W=2u
CS N2 0 1.3p
MP3 0 N2 N3 Vdd PMOS L=0.7u W=10u
MP4 N3 NRE Out Vdd PMOS L=0.7u W=10u

MC Out Out Vdd Vdd PMOS L=2u W=2u
CC Out 0 3p

*Testbench

.param Ipd_1 = 50p ! Photodiode current, range [50 pA, 750 pA]
.param VDD = 1.8 ! Supply voltage
.param EXPOSURETIME = 30m ! Exposure time, range [2 ms, 30 ms]

.param TRF = {EXPOSURETIME/100} ! Risetime and falltime of EXPOSURE and ERASE signals
.param PW = {EXPOSURETIME} ! Pulsewidth of EXPOSURE and ERASE signals
.param PERIOD = {EXPOSURETIME*10} ! Period for testbench sources
.param FS = 1k; ! Sampling clock frequency
.param CLK_PERIOD = {1/FS} ! Sampling clock period
.param EXPOSE_DLY = {CLK_PERIOD} ! Delay for EXPOSE signal
.param NRE_DLY = {2*CLK_PERIOD + EXPOSURETIME} ! Delay for NRE signal
.param ERASE_DLY = {6*CLK_PERIOD + EXPOSURETIME} ! Delay for ERASE signal

VDD Vdd 0 dc VDD
VEXPOSE Expose 0 dc 0 pulse(0 VDD EXPOSE_DLY TRF TRF EXPOSURETIME PERIOD)
VERASE Erase 0 dc 0 pulse(0 VDD ERASE_DLY TRF TRF CLK_PERIOD PERIOD)
VNRE NRE 0 dc 0 pulse(VDD 0 NRE_DLY TRF TRF CLK_PERIOD PERIOD)

.plot V(EXPOSE) V(ERASE) V(NRE) V(Out) V(N2) V(N3)
.plot V(out)

.subckt PhotoDiode  VDD N1_R1C1
I1_R1C1  VDD   N1_R1C1   DC  Ipd_1
d1 N1_R1C1 vdd dwell 1
.model dwell d cj0=1e-14 is=1e-12 m=0.5 bv=40
Cd1 N1_R1C1 VDD 30f
.ends 

[tran]
0.0001
0.060
X
X
0
[ana]
4 0
[end]
